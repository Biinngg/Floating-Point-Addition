library verilog;
use verilog.vl_types.all;
entity test_bench is
end test_bench;
